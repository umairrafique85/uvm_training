interface cuboid_inp_intf (input clk);

  logic [16-1:0] length;
  logic [16-1:0] width;
  logic [16-1:0] height;
  logic          valid ;

endinterface

 interface cuboid_out_intf (input clk);

  logic [32-1:0] area;
  logic [32-1:0] volm;
  logic          valid;

endinterface